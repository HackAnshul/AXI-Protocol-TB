package axi_test_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "axi_defines.sv"
 // `include "ram_env_pkg.sv"
  import axi_mas_agt_pkg::*;
  import axi_slv_agt_pkg::*;
  import axi_env_pkg::*;
  `include "axi_env_config.svh"

  `include "axi_base_test.sv"

  //testcases go below

endpackage
