`ifndef AXI_MAS_DEFINES_SV
`define AXI_MAS_DEFINES_SV

// `define ADDR_WIDTH 32 //MAS_ADDR
// `define DATA_WIDTH 32
// `define DRAIN_TIME 900000
// `define ID_X_WIDTH 8

`endif
