//HEADER
`ifndef AXI_DEFINES_SV
`define AXI_DEFINES_SV

`define ADDR_WIDTH 32
`define DATA_WIDTH 32
`define DRAIN_TIME 900000
`define ID_X_WIDTH 8

`endif
