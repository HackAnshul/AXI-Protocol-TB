`ifndef AXI_SLV_PKG_SV
`define AXI_SLV_PKG_SV
`include "axi_defines.svh"
  `include "axi_slv_inf.sv"
package axi_slv_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

`include "axi_slv_defines.sv"
  //`include "axi_slv_config.svh"

  import axi_mas_agt_pkg::*;
endpackage
`endif
