package axi_mas_agt_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "axi_defines.svh"
  `include "axi_mas_config.svh"
  `include "axi_mas_seq_item.sv"
  `include "axi_mas_seqr.sv"
  `include "axi_mas_drv.sv"
  `include "axi_mas_mon.sv"
  `include "axi_mas_agent.sv"

  `include "axi_mas_base_seqs.sv"
endpackage
