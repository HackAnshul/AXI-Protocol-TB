`ifndef AXI_SLV_DEFINES_SV
`define AXI_SLV_DEFINES_SV

// `define ADDR_WIDTH 32 //SLV_ADDR
// `define DATA_WIDTH 32
// `define DRAIN_TIME 900000
// `define ID_X_WIDTH 8

`endif
